`define FOO2 99

module foo2;
endmodule

module foo2_friend;
endmodule
