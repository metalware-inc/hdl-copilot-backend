`define ABC 2
