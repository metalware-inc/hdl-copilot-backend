module bad;
endmodule
fewf
