module m;
    initial begin
        $display("FOO: %d", `FOO);
    end
endmodule
