module main_tb;
    foo2 f2();

    foo2_foe f2f();
    foo1 f1();

    initial begin
        $display("FOO2: %d", `FOO2);
    end
endmodule
