`define FOO2 98

module foo2;
endmodule

module foo2_foe;
endmodule
