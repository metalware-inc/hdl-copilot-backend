`define FOO 3