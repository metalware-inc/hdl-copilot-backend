module foo (input logic rst, input logic clk);
endmodule