module foo_tb;
    wire clk, rst;
    foo f(clk, rst);
endmodule

