`define FOO1 2

module foo1;
endmodule
