module good;
endmodule
