`define WIDTH 4
